LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
-------------------------------------
ENTITY BinUnivCont IS
	GENERIC(N		  : INTEGER := 3;
			  MAX_COUNT: INTEGER := 5);
	PORT 	 (clk		  : IN	STD_LOGIC;
			  rst		  : IN	STD_LOGIC;
			  ena 	  : IN	STD_LOGIC;
			  syn_clr  : IN	STD_LOGIC;
			  load     : IN	STD_LOGIC;
			  up		  : IN	STD_LOGIC;
			  d 		  : IN	STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			  max_tick : OUT 	STD_LOGIC;
			  min_tick : OUT 	STD_LOGIC;
			  counter  : OUT	STD_LOGIC_VECTOR(N-1 DOWNTO 0)
			  );
END ENTITY BinUnivCont;
-------------------------------------
ARCHITECTURE rtl OF BinUnivCont IS
	--CONSTANT ONES 		:	UNSIGNED(N-1 DOWNTO 0) := (OTHERS => '1');
	CONSTANT ZEROS		:	UNSIGNED(N-1 DOWNTO 0) := (OTHERS => '0');
	
	SIGNAL count_s		: 	UNSIGNED(N-1 DOWNTO 0);
	SIGNAL count_next	: 	UNSIGNED(N-1 DOWNTO 0);
	SIGNAL max_reach  :  STD_LOGIC;
	SIGNAL min_reach  :  STD_LOGIC;
	SIGNAL max_up  	:  STD_LOGIC;
	SIGNAL min_up  	:  STD_LOGIC;
	
BEGIN

	-- NEXT STATE LOGIC
	count_next 	<= (OTHERS => '0')  		 WHEN ((syn_clr = '1') OR (max_up = '1'))	ELSE
						(TO_UNSIGNED(MAX_COUNT, N)) WHEN (min_up = '1')						ELSE
						UNSIGNED(d)	 	  		 WHEN load = '1'					  				ELSE
						count_s + 1		   	 WHEN (ena = '1' AND up = '1') 			 	ELSE
						count_s - 1	  	  		 WHEN (ena = '1' AND up = '0')  				ELSE
						count_s;
						 
	PROCESS(clk, rst)
		VARIABLE temp : UNSIGNED(N-1 DOWNTO 0);
	BEGIN
		IF(rst = '1') THEN
			temp := (OTHERS => '0');
		ELSIF (rising_edge(clk)) THEN
			IF (ena = '1') THEN 
				IF(temp <= TO_UNSIGNED(MAX_COUNT,N)) THEN
					temp := count_next;
				END IF;
			END IF;
		END IF;
		counter <= STD_LOGIC_VECTOR(temp);
		count_s <= temp;
	END PROCESS;
	-- OUTPUT LOGIC
	max_reach  <= '1' WHEN count_s = TO_UNSIGNED(MAX_COUNT,N)	ELSE '0';
	max_tick   <= max_reach;
	max_up     <= '1' WHEN (max_reach = '1' AND up = '1') ELSE '0';
	
	min_reach  <= '1' WHEN count_s = ZEROS	ELSE '0';	
	min_tick   <= min_reach;
	min_up	  <= '1' WHEN (min_reach = '1' AND up = '0') ELSE '0';
	
END ARCHITECTURE;